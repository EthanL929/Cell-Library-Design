magic
tech tsmc180
timestamp 1670606464
<< nwell >>
rect 0 429 264 866
<< polysilicon >>
rect 39 774 48 785
rect 79 774 88 785
rect 119 774 128 785
rect 159 774 168 785
rect 39 628 48 725
rect 79 628 88 725
rect 39 258 48 603
rect 79 258 88 603
rect 119 591 128 725
rect 119 258 128 566
rect 159 554 168 725
rect 159 258 168 529
rect 39 220 48 231
rect 79 220 88 231
rect 119 219 128 231
rect 159 160 168 231
<< ndiffusion >>
rect 36 231 39 258
rect 48 231 79 258
rect 88 231 119 258
rect 128 231 159 258
rect 168 231 171 258
<< pdiffusion >>
rect 36 725 39 774
rect 48 725 51 774
rect 76 725 79 774
rect 88 725 91 774
rect 116 725 119 774
rect 128 725 131 774
rect 156 725 159 774
rect 168 725 171 774
<< pohmic >>
rect 0 7 173 32
rect 198 7 264 32
<< nohmic >>
rect 0 834 51 859
rect 76 834 133 859
rect 158 834 264 859
<< ntransistor >>
rect 39 231 48 258
rect 79 231 88 258
rect 119 231 128 258
rect 159 231 168 258
<< ptransistor >>
rect 39 725 48 774
rect 79 725 88 774
rect 119 725 128 774
rect 159 725 168 774
<< polycontact >>
rect 25 603 50 628
rect 65 603 90 628
rect 110 566 135 591
rect 154 529 179 554
<< ndiffcontact >>
rect 11 231 36 258
rect 171 231 196 258
<< pdiffcontact >>
rect 11 725 36 774
rect 51 725 76 774
rect 91 725 116 774
rect 131 725 156 774
rect 171 725 196 774
<< psubstratetap >>
rect 173 7 198 32
<< nsubstratetap >>
rect 51 834 76 859
rect 133 834 158 859
<< metal1 >>
rect 0 834 51 859
rect 76 834 133 859
rect 158 834 264 859
rect 57 774 69 834
rect 138 774 150 834
rect 19 657 31 725
rect 97 657 109 725
rect 179 657 191 725
rect 19 645 222 657
rect 0 434 264 446
rect 0 401 264 413
rect 0 377 264 389
rect 0 353 264 365
rect 0 329 264 341
rect 18 280 222 292
rect 18 258 30 280
rect 178 32 190 231
rect 0 7 173 32
rect 198 7 264 32
<< m2contact >>
rect 222 642 247 667
rect 23 603 25 628
rect 25 603 48 628
rect 62 603 65 628
rect 65 603 87 628
rect 124 566 135 591
rect 135 566 149 591
rect 163 529 179 554
rect 179 529 188 554
rect 222 274 247 301
<< metal2 >>
rect 33 628 47 866
rect 66 628 80 866
rect 33 0 47 603
rect 66 0 80 603
rect 132 591 146 866
rect 132 0 146 566
rect 165 554 179 866
rect 231 667 245 866
rect 165 0 179 529
rect 231 301 245 642
rect 231 0 245 274
<< labels >>
rlabel metal1 0 329 0 341 3 nReset
rlabel metal1 0 353 0 365 3 Clock
rlabel metal1 0 377 0 389 3 Test
rlabel metal1 0 401 0 413 3 Scan
rlabel metal1 0 434 0 446 3 ScanReturn
rlabel metal1 0 7 0 32 3 GND!
rlabel metal1 0 834 0 859 3 Vdd!
rlabel metal2 33 866 47 866 5 A
rlabel metal2 33 0 47 0 1 A
rlabel metal2 66 866 80 866 5 B
rlabel metal2 66 0 80 0 1 B
rlabel metal2 132 866 146 866 5 C
rlabel metal2 132 0 146 0 1 C
rlabel metal2 165 866 179 866 5 D
rlabel metal2 165 0 179 0 1 D
rlabel metal2 231 866 245 866 5 Y
rlabel metal2 231 0 245 0 1 Y
rlabel metal1 264 7 264 32 7 GND!
rlabel metal1 264 377 264 389 7 Test
rlabel metal1 264 353 264 365 7 Clock
rlabel metal1 264 329 264 341 7 nReset
rlabel metal1 264 401 264 413 7 Scan
rlabel metal1 264 434 264 446 7 ScanReturn
rlabel metal1 264 834 264 859 7 Vdd!
<< end >>
