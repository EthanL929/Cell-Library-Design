magic
tech tsmc180
timestamp 1670606464
<< nwell >>
rect 0 429 429 866
<< polysilicon >>
rect 57 807 66 818
rect 95 807 104 818
rect 57 542 66 758
rect 95 683 104 758
rect 135 683 144 818
rect 173 807 182 818
rect 211 807 220 818
rect 173 746 182 758
rect 173 683 182 725
rect 211 683 220 758
rect 249 716 258 818
rect 287 807 296 818
rect 327 807 336 818
rect 287 746 296 783
rect 249 683 258 695
rect 287 683 296 725
rect 327 716 336 783
rect 327 683 336 695
rect 57 311 66 521
rect 95 374 104 634
rect 135 598 144 634
rect 173 598 182 634
rect 211 598 220 634
rect 249 598 258 634
rect 135 513 144 549
rect 95 353 101 374
rect 57 231 66 290
rect 57 222 68 231
rect 59 210 68 222
rect 95 210 104 353
rect 135 317 144 492
rect 173 317 182 549
rect 211 350 220 549
rect 211 317 220 329
rect 249 317 258 549
rect 287 422 296 634
rect 327 422 336 634
rect 367 598 376 818
rect 367 479 376 549
rect 287 401 298 422
rect 287 317 296 401
rect 327 311 336 401
rect 59 170 68 183
rect 57 161 68 170
rect 57 48 66 161
rect 95 108 104 183
rect 135 141 144 290
rect 173 210 182 290
rect 211 210 220 290
rect 173 171 182 183
rect 135 108 144 120
rect 173 108 182 150
rect 211 108 220 183
rect 249 168 258 290
rect 287 204 296 290
rect 327 210 336 290
rect 249 108 258 144
rect 287 168 296 183
rect 327 168 336 183
rect 95 48 104 81
rect 135 48 144 81
rect 173 48 182 81
rect 211 48 220 81
rect 249 48 258 81
rect 287 48 296 144
rect 327 117 336 144
rect 367 117 376 458
rect 309 108 336 117
rect 349 108 376 117
rect 309 48 318 108
rect 349 93 358 108
rect 349 48 358 66
<< ndiffusion >>
rect 130 290 135 317
rect 144 290 173 317
rect 182 290 211 317
rect 220 290 223 317
rect 244 290 249 317
rect 258 290 287 317
rect 296 290 301 317
rect 56 183 59 210
rect 68 183 95 210
rect 104 183 109 210
rect 170 183 173 210
rect 182 183 211 210
rect 220 183 223 210
rect 322 183 327 210
rect 336 183 341 210
rect 92 81 95 108
rect 104 81 135 108
rect 144 81 173 108
rect 182 81 211 108
rect 220 81 223 108
rect 244 81 249 108
rect 258 81 261 108
rect 344 66 349 93
rect 358 66 361 93
<< pdiffusion >>
rect 54 758 57 807
rect 66 758 71 807
rect 92 758 95 807
rect 104 758 109 807
rect 170 758 173 807
rect 182 758 187 807
rect 208 758 211 807
rect 220 758 223 807
rect 92 634 95 683
rect 104 634 109 683
rect 130 634 135 683
rect 144 634 149 683
rect 170 634 173 683
rect 182 634 187 683
rect 208 634 211 683
rect 220 634 223 683
rect 244 634 249 683
rect 258 634 261 683
rect 282 634 287 683
rect 296 634 301 683
rect 322 634 327 683
rect 336 634 341 683
rect 130 549 135 598
rect 144 549 149 598
rect 170 549 173 598
rect 182 549 187 598
rect 208 549 211 598
rect 220 549 223 598
rect 244 549 249 598
rect 258 549 261 598
rect 362 549 367 598
rect 376 549 379 598
<< pohmic >>
rect 0 11 9 32
rect 30 11 429 32
rect 0 7 429 11
<< nohmic >>
rect 0 855 429 859
rect 0 834 9 855
rect 30 834 429 855
<< ntransistor >>
rect 135 290 144 317
rect 173 290 182 317
rect 211 290 220 317
rect 249 290 258 317
rect 287 290 296 317
rect 59 183 68 210
rect 95 183 104 210
rect 173 183 182 210
rect 211 183 220 210
rect 327 183 336 210
rect 95 81 104 108
rect 135 81 144 108
rect 173 81 182 108
rect 211 81 220 108
rect 249 81 258 108
rect 349 66 358 93
<< ptransistor >>
rect 57 758 66 807
rect 95 758 104 807
rect 173 758 182 807
rect 211 758 220 807
rect 95 634 104 683
rect 135 634 144 683
rect 173 634 182 683
rect 211 634 220 683
rect 249 634 258 683
rect 287 634 296 683
rect 327 634 336 683
rect 135 549 144 598
rect 173 549 182 598
rect 211 549 220 598
rect 249 549 258 598
rect 367 549 376 598
<< polycontact >>
rect 163 725 184 746
rect 287 783 311 807
rect 327 783 351 807
rect 279 725 300 746
rect 237 695 258 716
rect 315 695 336 716
rect 51 521 72 542
rect 123 492 144 513
rect 101 353 122 374
rect 51 290 72 311
rect 206 329 227 350
rect 367 458 388 479
rect 322 401 343 422
rect 327 290 348 311
rect 163 150 184 171
rect 129 120 150 141
rect 275 183 296 204
rect 234 144 258 168
rect 287 144 311 168
rect 327 144 351 168
<< ndiffcontact >>
rect 109 290 130 317
rect 223 290 244 317
rect 301 290 322 317
rect 35 183 56 210
rect 109 183 130 210
rect 149 183 170 210
rect 223 183 244 210
rect 301 183 322 210
rect 341 183 362 210
rect 71 81 92 108
rect 223 81 244 108
rect 261 81 282 108
rect 323 66 344 93
rect 361 66 382 93
<< pdiffcontact >>
rect 33 758 54 807
rect 71 758 92 807
rect 109 758 130 807
rect 149 758 170 807
rect 187 758 208 807
rect 223 758 244 807
rect 71 634 92 683
rect 109 634 130 683
rect 149 634 170 683
rect 187 634 208 683
rect 223 634 244 683
rect 261 634 282 683
rect 301 634 322 683
rect 341 634 362 683
rect 109 549 130 598
rect 149 549 170 598
rect 187 549 208 598
rect 223 549 244 598
rect 261 549 282 598
rect 341 549 362 598
rect 379 549 400 598
<< psubstratetap >>
rect 9 11 30 32
<< nsubstratetap >>
rect 9 834 30 855
<< metal1 >>
rect 0 855 429 859
rect 0 834 9 855
rect 30 834 429 855
rect 33 807 45 834
rect 114 807 126 834
rect 154 807 166 834
rect 228 807 240 834
rect 33 622 45 758
rect 75 740 87 758
rect 75 728 163 740
rect 196 740 208 758
rect 196 728 279 740
rect 300 728 362 740
rect 114 701 237 713
rect 114 683 126 701
rect 192 683 204 701
rect 270 701 315 713
rect 270 683 282 701
rect 350 683 362 728
rect 75 622 87 634
rect 154 622 166 634
rect 227 622 239 634
rect 305 622 317 634
rect 33 610 395 622
rect 154 598 166 610
rect 227 598 239 610
rect 383 598 395 610
rect 282 586 341 598
rect 114 537 126 549
rect 192 537 204 549
rect 72 525 204 537
rect 266 509 278 549
rect 144 497 278 509
rect 0 470 80 482
rect 68 458 367 470
rect 0 434 429 446
rect 53 413 299 422
rect 0 410 322 413
rect 0 401 65 410
rect 287 401 322 410
rect 343 401 429 413
rect 77 389 275 398
rect 0 386 429 389
rect 0 377 89 386
rect 263 377 429 386
rect 0 353 101 365
rect 122 365 251 374
rect 122 362 429 365
rect 239 353 429 362
rect 0 329 206 341
rect 227 329 429 341
rect 72 290 109 302
rect 322 290 327 311
rect 227 256 239 290
rect 35 244 239 256
rect 35 210 47 244
rect 149 210 161 244
rect 251 234 357 246
rect 251 222 263 234
rect 232 210 263 222
rect 345 210 357 234
rect 296 183 301 204
rect 35 32 47 183
rect 118 171 130 183
rect 118 159 163 171
rect 150 120 382 132
rect 76 108 88 120
rect 370 93 382 120
rect 282 81 323 93
rect 228 32 240 81
rect 0 11 9 32
rect 30 11 429 32
rect 0 7 429 11
<< m2contact >>
rect 287 783 311 807
rect 327 783 351 807
rect 234 144 258 168
rect 287 144 311 168
rect 327 144 351 168
rect 70 120 94 144
<< metal2 >>
rect 297 807 311 866
rect 330 807 344 866
rect 297 168 311 783
rect 330 168 344 783
rect 94 130 258 144
rect 297 0 311 144
rect 330 0 344 144
<< labels >>
rlabel metal1 0 834 0 859 3 Vdd!
rlabel metal1 0 329 0 341 3 nReset
rlabel metal1 0 353 0 365 3 Clock
rlabel metal1 0 377 0 389 3 Test
rlabel metal1 0 401 0 413 3 Q
rlabel metal1 0 434 0 446 3 ScanReturn
rlabel metal1 0 470 0 482 3 nD
rlabel metal1 0 7 0 32 3 GND!
rlabel metal1 429 434 429 446 7 ScanReturn
rlabel metal1 429 353 429 365 7 Clock
rlabel metal1 429 377 429 389 7 Test
rlabel metal1 429 401 429 413 7 Q
rlabel metal1 429 329 429 341 7 nReset
rlabel metal1 429 834 429 859 7 Vdd!
rlabel metal1 429 7 429 32 7 GND!
rlabel metal2 297 0 311 0 1 nQ
rlabel metal2 330 0 344 0 1 Q
rlabel metal2 297 866 311 866 5 nQ
rlabel metal2 330 866 344 866 5 Q
<< end >>
