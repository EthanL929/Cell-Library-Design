magic
tech tsmc180
timestamp 1670606464
<< nwell >>
rect 0 429 594 866
<< polysilicon >>
rect 132 806 141 820
rect 198 806 207 812
rect 66 717 75 759
rect 331 779 340 796
rect 132 717 141 757
rect 198 717 207 757
rect 331 770 372 779
rect 264 717 273 753
rect 363 717 372 770
rect 462 717 471 757
rect 528 717 537 757
rect 66 426 75 668
rect 132 403 141 668
rect 66 155 75 401
rect 132 196 141 377
rect 198 194 207 668
rect 132 155 141 169
rect 198 155 207 170
rect 264 155 273 668
rect 363 629 372 668
rect 462 629 471 668
rect 363 195 372 580
rect 334 186 372 195
rect 334 155 343 163
rect 462 156 471 580
rect 528 428 537 668
rect 528 156 537 401
rect 66 59 75 128
rect 132 61 141 128
rect 198 63 207 128
rect 264 86 273 128
rect 334 88 343 128
rect 462 86 471 129
rect 528 65 537 129
rect 334 45 343 61
<< ndiffusion >>
rect 116 169 132 196
rect 141 169 146 196
rect 61 128 66 155
rect 75 128 132 155
rect 141 128 156 155
rect 177 128 198 155
rect 207 128 227 155
rect 250 128 264 155
rect 273 128 334 155
rect 343 128 386 155
rect 449 129 462 156
rect 471 129 528 156
rect 537 129 541 156
rect 328 61 334 88
rect 343 61 352 88
<< pdiffusion >>
rect 115 757 132 806
rect 141 757 160 806
rect 60 668 66 717
rect 75 668 93 717
rect 114 668 132 717
rect 141 668 161 717
rect 182 668 198 717
rect 207 668 226 717
rect 247 668 264 717
rect 273 668 323 717
rect 344 668 363 717
rect 372 668 381 717
rect 449 668 462 717
rect 471 668 490 717
rect 511 668 528 717
rect 537 668 541 717
rect 351 580 363 629
rect 372 580 387 629
<< pohmic >>
rect 0 30 594 32
rect 0 9 86 30
rect 107 9 157 30
rect 178 9 386 30
rect 409 9 456 30
rect 479 9 594 30
rect 0 7 594 9
<< nohmic >>
rect 0 858 594 859
rect 0 837 83 858
rect 104 837 155 858
rect 176 857 471 858
rect 176 837 406 857
rect 0 836 406 837
rect 429 837 471 857
rect 494 837 594 858
rect 429 836 594 837
rect 0 834 594 836
<< ntransistor >>
rect 132 169 141 196
rect 66 128 75 155
rect 132 128 141 155
rect 198 128 207 155
rect 264 128 273 155
rect 334 128 343 155
rect 462 129 471 156
rect 528 129 537 156
rect 334 61 343 88
<< ptransistor >>
rect 132 757 141 806
rect 66 668 75 717
rect 132 668 141 717
rect 198 668 207 717
rect 264 668 273 717
rect 363 668 372 717
rect 462 668 471 717
rect 528 668 537 717
rect 363 580 372 629
<< polycontact >>
rect 192 757 213 806
rect 326 796 349 820
rect 259 753 280 778
rect 60 401 81 426
rect 126 377 147 403
rect 191 170 213 194
rect 455 580 476 629
rect 321 163 344 186
rect 519 401 545 428
rect 256 65 281 86
rect 456 61 480 86
<< ndiffcontact >>
rect 95 169 116 196
rect 146 169 167 196
rect 40 128 61 155
rect 156 128 177 155
rect 227 128 250 155
rect 386 128 407 155
rect 428 129 449 156
rect 541 129 562 156
rect 307 61 328 88
rect 352 61 373 88
<< pdiffcontact >>
rect 94 757 115 806
rect 160 757 181 806
rect 39 668 60 717
rect 93 668 114 717
rect 161 668 182 717
rect 226 668 247 717
rect 323 668 344 717
rect 381 668 402 717
rect 428 668 449 717
rect 490 668 511 717
rect 541 668 562 717
rect 330 580 351 629
rect 387 580 408 629
<< psubstratetap >>
rect 86 9 107 30
rect 157 9 178 30
rect 386 9 409 30
rect 456 9 479 30
<< nsubstratetap >>
rect 83 837 104 858
rect 155 837 176 858
rect 406 836 429 857
rect 471 837 494 858
<< metal1 >>
rect 0 858 594 859
rect 0 837 83 858
rect 104 837 155 858
rect 176 857 471 858
rect 176 837 406 857
rect 0 836 406 837
rect 429 837 471 857
rect 494 837 594 858
rect 429 836 594 837
rect 0 834 594 836
rect 99 806 111 834
rect 181 757 192 806
rect 43 733 177 745
rect 43 717 55 733
rect 165 717 177 733
rect 230 717 242 834
rect 165 568 177 668
rect 299 608 311 834
rect 385 717 397 834
rect 433 737 557 749
rect 433 717 445 737
rect 545 717 557 737
rect 327 655 339 668
rect 495 655 507 668
rect 327 643 507 655
rect 299 596 330 608
rect 408 595 455 607
rect 545 568 557 668
rect 165 556 557 568
rect 177 499 567 511
rect 555 482 567 499
rect 555 470 594 482
rect 30 458 167 468
rect 30 456 572 458
rect 30 446 42 456
rect 155 446 572 456
rect 0 434 42 446
rect 560 434 594 446
rect 0 401 60 413
rect 0 377 126 389
rect 545 401 594 413
rect 147 377 594 389
rect 0 353 594 365
rect 0 329 594 341
rect 96 220 108 232
rect 47 208 444 220
rect 47 155 59 208
rect 167 170 191 194
rect 99 32 111 169
rect 391 155 403 208
rect 432 156 444 208
rect 161 32 173 128
rect 231 115 243 128
rect 544 115 556 129
rect 231 103 556 115
rect 373 67 456 79
rect 311 32 323 61
rect 0 30 594 32
rect 0 9 86 30
rect 107 9 157 30
rect 178 9 386 30
rect 409 9 456 30
rect 479 9 594 30
rect 0 7 594 9
<< m2contact >>
rect 259 753 280 778
rect 93 676 114 700
rect 326 796 349 820
rect 154 493 177 516
rect 90 232 116 260
rect 321 163 344 186
rect 256 65 281 86
<< metal2 >>
rect 264 778 278 866
rect 330 820 344 866
rect 96 514 110 676
rect 96 500 154 514
rect 96 260 110 500
rect 264 0 278 65
rect 330 0 344 163
<< labels >>
rlabel metal2 330 0 344 0 1 Load
rlabel metal2 264 0 278 0 1 D
rlabel metal1 0 7 0 32 3 GND!
rlabel metal1 0 377 0 389 3 Test
rlabel metal1 0 353 0 365 3 Clock
rlabel metal1 0 329 0 341 3 nReset
rlabel metal1 0 401 0 413 3 SDI
rlabel metal1 0 434 0 446 3 ScanReturn
rlabel metal1 594 7 594 32 7 GND!
rlabel metal1 594 353 594 365 7 Clock
rlabel metal1 594 377 594 389 7 Test
rlabel metal1 594 329 594 341 7 nReset
rlabel metal1 594 401 594 413 7 Q
rlabel metal1 594 434 594 446 7 ScanReturn
rlabel metal1 594 470 594 482 7 nD
rlabel metal1 0 834 0 859 3 Vdd!
rlabel metal2 264 866 278 866 5 D
rlabel metal2 330 866 344 866 5 Load
rlabel metal1 594 834 594 859 7 Vdd!
<< end >>
