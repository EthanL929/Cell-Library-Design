magic
tech tsmc180
timestamp 1670606464
<< nwell >>
rect 250 429 1650 866
<< polysilicon >>
rect 330 805 339 816
rect 414 805 423 816
rect 485 805 494 816
rect 557 805 566 816
rect 593 805 602 816
rect 664 805 673 816
rect 701 805 710 816
rect 737 805 746 816
rect 810 805 819 816
rect 330 420 339 756
rect 330 93 339 395
rect 414 119 423 749
rect 485 206 494 654
rect 557 399 566 601
rect 593 399 602 601
rect 881 803 890 814
rect 963 804 972 815
rect 999 804 1008 815
rect 557 390 602 399
rect 485 116 494 181
rect 557 176 566 390
rect 557 136 566 151
rect 593 136 602 390
rect 664 347 673 431
rect 701 347 710 431
rect 737 347 746 431
rect 664 338 746 347
rect 664 238 673 338
rect 664 201 673 213
rect 701 201 710 338
rect 737 201 746 338
rect 414 80 423 94
rect 330 54 339 66
rect 810 119 819 749
rect 881 211 890 652
rect 1070 803 1079 814
rect 1107 803 1116 814
rect 1143 803 1152 815
rect 1239 806 1248 817
rect 963 398 972 600
rect 999 398 1008 600
rect 1310 804 1319 815
rect 1392 805 1401 816
rect 1428 805 1437 816
rect 1499 805 1508 816
rect 1536 805 1545 816
rect 1572 805 1581 816
rect 963 389 1008 398
rect 881 116 890 186
rect 963 175 972 389
rect 963 136 972 150
rect 999 136 1008 389
rect 1070 345 1079 429
rect 1107 345 1116 429
rect 1143 345 1152 429
rect 1070 336 1152 345
rect 1070 236 1079 336
rect 1070 199 1079 211
rect 1107 199 1116 336
rect 1143 199 1152 336
rect 810 80 819 94
rect 414 48 423 59
rect 485 47 494 59
rect 557 48 566 59
rect 593 48 602 59
rect 664 50 673 61
rect 701 50 710 61
rect 737 50 746 61
rect 1239 121 1248 750
rect 1310 210 1319 653
rect 1392 399 1401 601
rect 1428 399 1437 601
rect 1392 390 1437 399
rect 1310 116 1319 185
rect 1392 174 1401 390
rect 1392 136 1401 149
rect 1428 136 1437 390
rect 1499 346 1508 431
rect 1536 346 1545 431
rect 1572 346 1581 431
rect 1499 337 1581 346
rect 1499 236 1508 337
rect 1499 199 1508 211
rect 1536 199 1545 337
rect 1572 199 1581 337
rect 1239 82 1248 96
rect 810 48 819 59
rect 881 48 890 59
rect 963 48 972 59
rect 999 48 1008 59
rect 1070 48 1079 59
rect 1107 48 1116 59
rect 1143 48 1152 59
rect 1239 50 1248 61
rect 1310 48 1319 59
rect 1392 47 1401 59
rect 1428 47 1437 59
rect 1499 48 1508 59
rect 1536 48 1545 59
rect 1572 48 1581 59
<< ndiffusion >>
rect 327 66 330 93
rect 339 66 342 93
rect 411 59 414 80
rect 423 59 426 80
rect 482 59 485 116
rect 494 59 497 116
rect 554 59 557 136
rect 566 59 569 136
rect 590 59 593 136
rect 602 59 605 136
rect 661 61 664 201
rect 673 61 677 201
rect 698 61 701 201
rect 710 61 713 201
rect 734 61 737 201
rect 746 61 749 201
rect 807 59 810 80
rect 819 59 822 80
rect 878 59 881 116
rect 890 59 893 116
rect 960 59 963 136
rect 972 59 975 136
rect 996 59 999 136
rect 1008 59 1011 136
rect 1067 59 1070 199
rect 1079 59 1083 199
rect 1104 59 1107 199
rect 1116 59 1119 199
rect 1140 59 1143 199
rect 1152 59 1155 199
rect 1236 61 1239 82
rect 1248 61 1251 82
rect 1307 59 1310 116
rect 1319 59 1322 116
rect 1389 59 1392 136
rect 1401 59 1404 136
rect 1425 59 1428 136
rect 1437 59 1440 136
rect 1496 59 1499 199
rect 1508 59 1512 199
rect 1533 59 1536 199
rect 1545 59 1548 199
rect 1569 59 1572 199
rect 1581 59 1584 199
<< pdiffusion >>
rect 327 756 330 805
rect 339 756 342 805
rect 411 749 414 805
rect 423 749 426 805
rect 482 654 485 805
rect 494 654 497 805
rect 554 601 557 805
rect 566 601 569 805
rect 590 601 593 805
rect 602 601 605 805
rect 661 431 664 805
rect 673 431 677 805
rect 698 431 701 805
rect 710 431 713 805
rect 734 431 737 805
rect 746 431 749 805
rect 807 749 810 805
rect 819 749 822 805
rect 878 652 881 803
rect 890 652 893 803
rect 960 600 963 804
rect 972 600 975 804
rect 996 600 999 804
rect 1008 600 1011 804
rect 1067 429 1070 803
rect 1079 429 1083 803
rect 1104 429 1107 803
rect 1116 429 1119 803
rect 1140 429 1143 803
rect 1152 429 1155 803
rect 1236 750 1239 806
rect 1248 750 1251 806
rect 1307 653 1310 804
rect 1319 653 1322 804
rect 1389 601 1392 805
rect 1401 601 1404 805
rect 1425 601 1428 805
rect 1437 601 1440 805
rect 1496 431 1499 805
rect 1508 431 1512 805
rect 1533 431 1536 805
rect 1545 431 1548 805
rect 1569 431 1572 805
rect 1581 431 1584 805
<< pohmic >>
rect 260 31 1650 32
rect 260 9 333 31
rect 356 30 1650 31
rect 356 29 1486 30
rect 356 9 666 29
rect 260 7 666 9
rect 689 7 1066 29
rect 1089 8 1486 29
rect 1509 8 1650 30
rect 1089 7 1650 8
<< nohmic >>
rect 250 857 630 859
rect 250 835 329 857
rect 352 837 630 857
rect 653 858 1650 859
rect 653 837 1030 858
rect 352 836 1030 837
rect 1053 836 1458 858
rect 1481 836 1650 858
rect 352 835 1650 836
rect 250 834 1650 835
<< ntransistor >>
rect 330 66 339 93
rect 414 59 423 80
rect 485 59 494 116
rect 557 59 566 136
rect 593 59 602 136
rect 664 61 673 201
rect 701 61 710 201
rect 737 61 746 201
rect 810 59 819 80
rect 881 59 890 116
rect 963 59 972 136
rect 999 59 1008 136
rect 1070 59 1079 199
rect 1107 59 1116 199
rect 1143 59 1152 199
rect 1239 61 1248 82
rect 1310 59 1319 116
rect 1392 59 1401 136
rect 1428 59 1437 136
rect 1499 59 1508 199
rect 1536 59 1545 199
rect 1572 59 1581 199
<< ptransistor >>
rect 330 756 339 805
rect 414 749 423 805
rect 485 654 494 805
rect 557 601 566 805
rect 593 601 602 805
rect 664 431 673 805
rect 701 431 710 805
rect 737 431 746 805
rect 810 749 819 805
rect 881 652 890 803
rect 963 600 972 804
rect 999 600 1008 804
rect 1070 429 1079 803
rect 1107 429 1116 803
rect 1143 429 1152 803
rect 1239 750 1248 806
rect 1310 653 1319 804
rect 1392 601 1401 805
rect 1428 601 1437 805
rect 1499 431 1508 805
rect 1536 431 1545 805
rect 1572 431 1581 805
<< polycontact >>
rect 320 395 345 420
rect 474 181 499 206
rect 402 94 427 119
rect 547 151 572 176
rect 654 213 679 238
rect 872 186 897 211
rect 799 94 824 119
rect 953 150 978 175
rect 1060 211 1085 236
rect 1302 185 1327 210
rect 1228 96 1253 121
rect 1382 149 1407 174
rect 1490 211 1515 236
<< ndiffcontact >>
rect 306 66 327 93
rect 342 66 363 93
rect 390 59 411 80
rect 426 59 447 80
rect 461 59 482 116
rect 497 59 518 116
rect 533 59 554 136
rect 569 59 590 136
rect 605 59 626 136
rect 640 61 661 201
rect 677 61 698 201
rect 713 61 734 201
rect 749 61 770 201
rect 786 59 807 80
rect 822 59 843 80
rect 857 59 878 116
rect 893 59 914 116
rect 939 59 960 136
rect 975 59 996 136
rect 1011 59 1032 136
rect 1046 59 1067 199
rect 1083 59 1104 199
rect 1119 59 1140 199
rect 1155 59 1176 199
rect 1215 61 1236 82
rect 1251 61 1272 82
rect 1286 59 1307 116
rect 1322 59 1343 116
rect 1368 59 1389 136
rect 1404 59 1425 136
rect 1440 59 1461 136
rect 1475 59 1496 199
rect 1512 59 1533 199
rect 1548 59 1569 199
rect 1584 59 1605 199
<< pdiffcontact >>
rect 306 756 327 805
rect 342 756 363 805
rect 390 749 411 805
rect 426 749 447 805
rect 461 654 482 805
rect 497 654 518 805
rect 533 601 554 805
rect 569 601 590 805
rect 605 601 626 805
rect 640 431 661 805
rect 677 431 698 805
rect 713 431 734 805
rect 749 431 770 805
rect 786 749 807 805
rect 822 749 843 805
rect 857 652 878 803
rect 893 652 914 803
rect 939 600 960 804
rect 975 600 996 804
rect 1011 600 1032 804
rect 1046 429 1067 803
rect 1083 429 1104 803
rect 1119 429 1140 803
rect 1155 429 1176 803
rect 1215 750 1236 806
rect 1251 750 1272 806
rect 1286 653 1307 804
rect 1322 653 1343 804
rect 1368 601 1389 805
rect 1404 601 1425 805
rect 1440 601 1461 805
rect 1475 431 1496 805
rect 1512 431 1533 805
rect 1548 431 1569 805
rect 1584 431 1605 805
<< psubstratetap >>
rect 333 9 356 31
rect 666 7 689 29
rect 1066 7 1089 29
rect 1486 8 1509 30
<< nsubstratetap >>
rect 329 835 352 857
rect 630 837 653 859
rect 1030 836 1053 858
rect 1458 836 1481 858
<< metal1 >>
rect 250 857 630 859
rect 250 835 329 857
rect 352 837 630 857
rect 653 858 1650 859
rect 653 837 1030 858
rect 352 836 1030 837
rect 1053 836 1458 858
rect 1481 836 1650 858
rect 352 835 1650 836
rect 250 834 1650 835
rect 307 805 320 834
rect 394 805 407 834
rect 465 805 478 834
rect 537 805 550 834
rect 609 805 622 834
rect 645 805 658 834
rect 718 805 731 834
rect 790 805 803 834
rect 861 803 874 834
rect 944 804 957 834
rect 1015 804 1028 834
rect 1052 803 1065 834
rect 1123 803 1136 834
rect 1219 806 1232 834
rect 1290 804 1303 834
rect 1372 805 1385 834
rect 1445 805 1458 834
rect 1479 805 1492 834
rect 1552 805 1565 834
rect 1618 446 1630 680
rect 1618 434 1650 446
rect 345 401 1447 413
rect 1486 401 1650 413
rect 1486 323 1498 401
rect 1535 377 1650 389
rect 289 311 1498 323
rect 1582 353 1650 365
rect 1582 292 1594 353
rect 1180 280 1594 292
rect 1606 329 1650 341
rect 1606 260 1618 329
rect 772 248 1618 260
rect 592 219 654 231
rect 449 187 474 199
rect 520 152 547 164
rect 311 32 324 66
rect 394 32 407 59
rect 845 195 872 207
rect 998 217 1060 229
rect 917 157 953 169
rect 461 32 474 59
rect 538 32 551 59
rect 610 32 623 59
rect 643 32 656 61
rect 717 32 730 61
rect 790 32 803 59
rect 1274 193 1302 205
rect 1427 217 1490 229
rect 1346 155 1382 167
rect 1219 82 1232 84
rect 857 32 870 59
rect 941 32 954 59
rect 1014 32 1027 59
rect 1050 32 1063 59
rect 1122 32 1135 59
rect 1219 32 1232 61
rect 1286 32 1299 59
rect 1372 32 1385 59
rect 1443 32 1456 59
rect 1479 32 1492 59
rect 1552 32 1565 59
rect 260 31 1650 32
rect 260 9 333 31
rect 356 30 1650 31
rect 356 29 1486 30
rect 356 9 666 29
rect 260 7 666 9
rect 689 7 1066 29
rect 1089 8 1486 29
rect 1509 8 1650 30
rect 1089 7 1650 8
<< m2contact >>
rect 31 834 250 859
rect 343 756 362 803
rect 428 749 447 805
rect 499 654 518 805
rect 570 601 589 805
rect 678 431 697 805
rect 750 431 769 805
rect 824 749 843 805
rect 895 652 914 803
rect 976 600 995 804
rect 1084 429 1103 803
rect 1156 429 1175 803
rect 1253 750 1272 806
rect 1324 653 1343 804
rect 1405 601 1424 805
rect 1513 431 1532 805
rect 1585 431 1604 805
rect 1618 680 1643 705
rect 1447 394 1472 419
rect 264 299 289 324
rect 1510 364 1535 389
rect 1155 272 1180 297
rect 747 241 772 266
rect 567 209 592 234
rect 424 174 449 199
rect 495 142 520 167
rect 390 94 402 119
rect 402 94 415 119
rect 342 66 363 93
rect 426 59 447 80
rect 447 59 449 80
rect 426 56 449 59
rect 499 59 518 116
rect 570 59 589 136
rect 678 61 697 201
rect 750 61 769 201
rect 820 182 845 207
rect 973 207 998 232
rect 892 147 917 172
rect 786 94 799 119
rect 799 94 811 119
rect 822 59 843 80
rect 822 55 843 59
rect 895 59 914 116
rect 976 59 995 136
rect 1084 59 1103 199
rect 1156 59 1175 199
rect 1249 180 1274 205
rect 1402 207 1427 232
rect 1321 145 1346 170
rect 1215 96 1228 121
rect 1228 96 1240 121
rect 1251 61 1272 82
rect 1251 57 1272 61
rect 1324 59 1343 116
rect 1405 59 1424 136
rect 1513 59 1532 199
rect 1585 59 1604 199
<< metal2 >>
rect 0 859 250 866
rect 0 834 31 859
rect 0 0 250 834
rect 264 724 278 866
rect 347 724 361 756
rect 264 710 361 724
rect 264 0 278 299
rect 347 93 361 710
rect 396 119 410 866
rect 429 199 443 749
rect 396 0 410 94
rect 429 80 443 174
rect 502 167 516 654
rect 573 234 587 601
rect 681 408 695 431
rect 753 408 767 431
rect 681 394 767 408
rect 502 116 516 142
rect 573 136 587 209
rect 681 201 695 394
rect 753 266 767 394
rect 753 201 767 241
rect 792 119 806 866
rect 825 207 839 749
rect 898 186 912 652
rect 979 232 993 600
rect 1087 404 1101 429
rect 1159 404 1173 429
rect 1087 390 1173 404
rect 792 0 806 94
rect 825 80 839 182
rect 898 172 913 186
rect 898 146 913 147
rect 898 116 912 146
rect 979 136 993 207
rect 1087 199 1101 390
rect 1159 297 1173 390
rect 1159 199 1173 272
rect 1221 121 1235 866
rect 1458 819 1632 833
rect 1254 205 1268 750
rect 1221 0 1235 96
rect 1254 82 1268 180
rect 1327 170 1341 653
rect 1408 232 1422 601
rect 1458 419 1472 819
rect 1618 705 1632 819
rect 1516 405 1530 431
rect 1588 405 1602 431
rect 1516 389 1602 405
rect 1535 388 1602 389
rect 1327 116 1341 145
rect 1408 136 1422 207
rect 1516 199 1530 364
rect 1588 199 1602 388
<< labels >>
rlabel metal1 1650 329 1650 341 7 nResetOut
rlabel metal1 1650 353 1650 365 7 ClockOut
rlabel metal1 1650 377 1650 389 7 TestOut
rlabel metal1 1650 401 1650 413 7 SDI
rlabel metal1 1650 434 1650 446 7 nSDO
rlabel metal1 1650 834 1650 859 7 Vdd!
rlabel metal1 1650 7 1650 32 7 GND!
rlabel metal2 264 0 278 0 1 SDI
rlabel metal2 396 0 410 0 1 nReset
rlabel metal2 792 0 806 0 1 Clock
rlabel metal2 1221 0 1235 0 1 Test
rlabel metal2 1221 866 1235 866 5 Test
rlabel metal2 792 866 806 866 5 Clock
rlabel metal2 396 866 410 866 5 nReset
rlabel metal2 264 866 278 866 5 SDO
rlabel metal2 0 866 250 866 5 Vdd!
rlabel metal2 0 0 250 0 1 Vdd!
<< end >>
