magic
tech tsmc180
timestamp 1670623449
<< nwell >>
rect 0 429 759 866
<< polysilicon >>
rect 66 717 75 811
rect 132 806 141 818
rect 198 806 207 818
rect 387 807 396 818
rect 425 807 434 818
rect 132 717 141 757
rect 198 717 207 757
rect 264 717 273 769
rect 66 434 75 668
rect 66 127 75 409
rect 132 399 141 668
rect 132 127 141 377
rect 198 127 207 668
rect 264 214 273 668
rect 387 542 396 758
rect 425 683 434 758
rect 465 683 474 818
rect 503 807 512 818
rect 541 807 550 818
rect 503 746 512 758
rect 503 683 512 725
rect 541 683 550 758
rect 579 716 588 818
rect 617 807 626 818
rect 657 807 666 818
rect 617 746 626 783
rect 579 683 588 695
rect 617 683 626 725
rect 657 716 666 783
rect 657 683 666 695
rect 387 311 396 521
rect 425 374 434 634
rect 465 598 474 634
rect 503 598 512 634
rect 541 598 550 634
rect 579 598 588 634
rect 465 513 474 549
rect 425 353 431 374
rect 387 231 396 290
rect 387 222 398 231
rect 389 210 398 222
rect 425 210 434 353
rect 465 317 474 492
rect 503 317 512 549
rect 541 350 550 549
rect 541 317 550 329
rect 579 317 588 549
rect 617 422 626 634
rect 657 422 666 634
rect 697 598 706 818
rect 697 479 706 549
rect 617 401 628 422
rect 617 317 626 401
rect 657 311 666 401
rect 264 127 273 189
rect 389 170 398 183
rect 387 161 398 170
rect 66 37 75 100
rect 132 86 141 100
rect 198 86 207 100
rect 264 85 273 100
rect 132 38 141 59
rect 198 37 207 59
rect 387 48 396 161
rect 425 108 434 183
rect 465 141 474 290
rect 503 210 512 290
rect 541 210 550 290
rect 503 171 512 183
rect 465 108 474 120
rect 503 108 512 150
rect 541 108 550 183
rect 579 168 588 290
rect 617 204 626 290
rect 657 210 666 290
rect 579 108 588 144
rect 617 168 626 183
rect 657 168 666 183
rect 425 48 434 81
rect 465 48 474 81
rect 503 48 512 81
rect 541 48 550 81
rect 579 48 588 81
rect 617 48 626 144
rect 657 117 666 144
rect 697 117 706 458
rect 639 108 666 117
rect 679 108 706 117
rect 639 48 648 108
rect 679 93 688 108
rect 679 48 688 66
<< ndiffusion >>
rect 460 290 465 317
rect 474 290 503 317
rect 512 290 541 317
rect 550 290 553 317
rect 574 290 579 317
rect 588 290 617 317
rect 626 290 631 317
rect 386 183 389 210
rect 398 183 425 210
rect 434 183 439 210
rect 59 100 66 127
rect 75 100 132 127
rect 141 100 156 127
rect 177 100 198 127
rect 207 100 264 127
rect 273 100 283 127
rect 116 59 132 86
rect 141 59 155 86
rect 500 183 503 210
rect 512 183 541 210
rect 550 183 553 210
rect 652 183 657 210
rect 666 183 671 210
rect 422 81 425 108
rect 434 81 465 108
rect 474 81 503 108
rect 512 81 541 108
rect 550 81 553 108
rect 574 81 579 108
rect 588 81 591 108
rect 674 66 679 93
rect 688 66 691 93
<< pdiffusion >>
rect 115 757 132 806
rect 141 757 160 806
rect 384 758 387 807
rect 396 758 401 807
rect 422 758 425 807
rect 434 758 439 807
rect 61 668 66 717
rect 75 668 93 717
rect 114 690 132 717
rect 118 668 132 690
rect 141 668 161 717
rect 182 668 198 717
rect 207 668 226 717
rect 247 668 264 717
rect 273 668 282 717
rect 500 758 503 807
rect 512 758 517 807
rect 538 758 541 807
rect 550 758 553 807
rect 422 634 425 683
rect 434 634 439 683
rect 460 634 465 683
rect 474 634 479 683
rect 500 634 503 683
rect 512 634 517 683
rect 538 634 541 683
rect 550 634 553 683
rect 574 634 579 683
rect 588 634 591 683
rect 612 634 617 683
rect 626 634 631 683
rect 652 634 657 683
rect 666 634 671 683
rect 460 549 465 598
rect 474 549 479 598
rect 500 549 503 598
rect 512 549 517 598
rect 538 549 541 598
rect 550 549 553 598
rect 574 549 579 598
rect 588 549 591 598
rect 692 549 697 598
rect 706 549 709 598
<< pohmic >>
rect 0 30 339 32
rect 0 9 86 30
rect 107 9 157 30
rect 178 11 339 30
rect 360 11 759 32
rect 178 9 759 11
rect 0 7 759 9
<< nohmic >>
rect 0 837 83 859
rect 104 837 155 859
rect 176 855 759 859
rect 176 837 339 855
rect 0 834 339 837
rect 360 834 759 855
<< ntransistor >>
rect 465 290 474 317
rect 503 290 512 317
rect 541 290 550 317
rect 579 290 588 317
rect 617 290 626 317
rect 389 183 398 210
rect 425 183 434 210
rect 66 100 75 127
rect 132 100 141 127
rect 198 100 207 127
rect 264 100 273 127
rect 132 59 141 86
rect 503 183 512 210
rect 541 183 550 210
rect 657 183 666 210
rect 425 81 434 108
rect 465 81 474 108
rect 503 81 512 108
rect 541 81 550 108
rect 579 81 588 108
rect 679 66 688 93
<< ptransistor >>
rect 132 757 141 806
rect 387 758 396 807
rect 425 758 434 807
rect 66 668 75 717
rect 132 668 141 717
rect 198 668 207 717
rect 264 668 273 717
rect 503 758 512 807
rect 541 758 550 807
rect 425 634 434 683
rect 465 634 474 683
rect 503 634 512 683
rect 541 634 550 683
rect 579 634 588 683
rect 617 634 626 683
rect 657 634 666 683
rect 465 549 474 598
rect 503 549 512 598
rect 541 549 550 598
rect 579 549 588 598
rect 697 549 706 598
<< polycontact >>
rect 192 757 213 806
rect 57 409 82 434
rect 127 377 148 399
rect 493 725 514 746
rect 617 783 641 807
rect 657 783 681 807
rect 609 725 630 746
rect 567 695 588 716
rect 645 695 666 716
rect 381 521 402 542
rect 453 492 474 513
rect 431 353 452 374
rect 381 290 402 311
rect 260 189 285 214
rect 536 329 557 350
rect 697 458 718 479
rect 652 401 673 422
rect 657 290 678 311
rect 191 59 212 86
rect 493 150 514 171
rect 459 120 480 141
rect 605 183 626 204
rect 564 144 588 168
rect 617 144 641 168
rect 657 144 681 168
<< ndiffcontact >>
rect 439 290 460 317
rect 553 290 574 317
rect 631 290 652 317
rect 365 183 386 210
rect 439 183 460 210
rect 38 100 59 127
rect 156 100 177 127
rect 283 100 304 127
rect 95 59 116 86
rect 155 59 176 86
rect 479 183 500 210
rect 553 183 574 210
rect 631 183 652 210
rect 671 183 692 210
rect 401 81 422 108
rect 553 81 574 108
rect 591 81 612 108
rect 653 66 674 93
rect 691 66 712 93
<< pdiffcontact >>
rect 94 757 115 806
rect 160 757 181 806
rect 363 758 384 807
rect 401 758 422 807
rect 439 758 460 807
rect 40 668 61 717
rect 93 690 114 717
rect 93 665 118 690
rect 161 668 182 717
rect 226 668 247 717
rect 282 668 303 717
rect 479 758 500 807
rect 517 758 538 807
rect 553 758 574 807
rect 401 634 422 683
rect 439 634 460 683
rect 479 634 500 683
rect 517 634 538 683
rect 553 634 574 683
rect 591 634 612 683
rect 631 634 652 683
rect 671 634 692 683
rect 439 549 460 598
rect 479 549 500 598
rect 517 549 538 598
rect 553 549 574 598
rect 591 549 612 598
rect 671 549 692 598
rect 709 549 730 598
<< psubstratetap >>
rect 86 9 107 30
rect 157 9 178 30
rect 339 11 360 32
<< nsubstratetap >>
rect 83 837 104 858
rect 155 837 176 858
rect 339 834 360 855
<< metal1 >>
rect 0 858 759 859
rect 0 837 83 858
rect 104 837 155 858
rect 176 855 759 858
rect 176 837 339 855
rect 0 834 339 837
rect 360 834 759 855
rect 99 806 111 834
rect 181 757 192 806
rect 45 730 177 742
rect 45 717 57 730
rect 165 717 177 730
rect 231 717 243 834
rect 363 807 375 834
rect 444 807 456 834
rect 484 807 496 834
rect 558 807 570 834
rect 167 656 179 668
rect 286 656 298 668
rect 167 644 298 656
rect 363 622 375 758
rect 405 740 417 758
rect 405 728 493 740
rect 526 740 538 758
rect 526 728 609 740
rect 630 728 692 740
rect 444 701 567 713
rect 444 683 456 701
rect 522 683 534 701
rect 600 701 645 713
rect 600 683 612 701
rect 680 683 692 728
rect 405 622 417 634
rect 484 622 496 634
rect 557 622 569 634
rect 635 622 647 634
rect 363 610 725 622
rect 484 598 496 610
rect 557 598 569 610
rect 713 598 725 610
rect 612 586 671 598
rect 444 537 456 549
rect 522 537 534 549
rect 402 525 534 537
rect 596 509 608 549
rect 474 497 608 509
rect 179 482 312 490
rect 179 478 410 482
rect 300 470 410 478
rect 9 449 229 461
rect 398 458 697 470
rect 9 446 21 449
rect 0 434 21 446
rect 217 446 229 449
rect 217 434 759 446
rect 33 415 57 427
rect 33 413 45 415
rect 0 401 45 413
rect 383 413 629 422
rect 330 410 652 413
rect 330 401 395 410
rect 617 401 652 410
rect 673 401 759 413
rect 0 377 127 389
rect 407 389 605 398
rect 148 386 759 389
rect 148 377 419 386
rect 593 377 759 386
rect 0 353 431 365
rect 452 365 581 374
rect 452 362 759 365
rect 569 353 759 362
rect 0 329 536 341
rect 557 329 759 341
rect 402 290 439 302
rect 652 290 657 311
rect 557 256 569 290
rect 365 244 569 256
rect 365 210 377 244
rect 479 210 491 244
rect 581 234 687 246
rect 581 222 593 234
rect 562 210 593 222
rect 675 210 687 234
rect 626 183 631 204
rect 43 32 55 100
rect 176 59 191 86
rect 100 32 112 59
rect 288 32 300 100
rect 365 32 377 183
rect 448 171 460 183
rect 448 159 493 171
rect 480 120 712 132
rect 406 108 418 120
rect 700 93 712 120
rect 612 81 653 93
rect 558 32 570 81
rect 0 30 339 32
rect 0 9 86 30
rect 107 9 157 30
rect 178 11 339 30
rect 360 11 759 32
rect 178 9 759 11
rect 0 7 759 9
<< m2contact >>
rect 617 783 641 807
rect 657 783 681 807
rect 93 665 118 690
rect 154 473 179 498
rect 260 189 285 214
rect 156 100 177 127
rect 564 144 588 168
rect 617 144 641 168
rect 657 144 681 168
rect 400 120 424 144
<< metal2 >>
rect 95 493 109 665
rect 95 479 154 493
rect 159 127 173 473
rect 264 214 278 866
rect 627 807 641 866
rect 660 807 674 866
rect 264 0 278 189
rect 627 168 641 783
rect 660 168 674 783
rect 424 130 588 144
rect 627 0 641 144
rect 660 0 674 144
<< labels >>
rlabel metal2 264 866 278 866 5 D
rlabel metal1 0 834 0 859 3 Vdd!
rlabel metal1 0 434 0 446 3 ScanReturn
rlabel metal1 0 401 0 413 3 SDI
rlabel metal1 0 377 0 389 3 Test
rlabel metal1 0 353 0 365 3 Clock
rlabel metal1 0 329 0 341 3 nReset
rlabel metal1 0 7 0 32 3 GND!
rlabel metal1 759 434 759 446 7 ScanReturn
rlabel metal1 759 353 759 365 7 Clock
rlabel metal1 759 377 759 389 7 Test
rlabel metal1 759 401 759 413 7 Q
rlabel metal1 759 329 759 341 7 nReset
rlabel metal1 759 834 759 859 7 Vdd!
rlabel metal1 759 7 759 32 7 GND!
rlabel metal2 627 0 641 0 1 nQ
rlabel metal2 660 0 674 0 1 Q
rlabel metal2 627 866 641 866 5 nQ
rlabel metal2 660 866 674 866 5 Q
rlabel metal2 264 0 278 0 1 D
<< end >>
