magic
tech tsmc180
timestamp 1670623489
<< nwell >>
rect 0 429 1023 866
<< polysilicon >>
rect 132 806 141 820
rect 198 806 207 812
rect 66 717 75 759
rect 651 807 660 818
rect 689 807 698 818
rect 331 779 340 792
rect 132 717 141 757
rect 198 717 207 757
rect 331 770 372 779
rect 264 717 273 749
rect 363 717 372 770
rect 462 717 471 757
rect 528 717 537 757
rect 66 426 75 668
rect 132 401 141 668
rect 66 155 75 401
rect 132 196 141 377
rect 198 194 207 668
rect 132 155 141 169
rect 198 155 207 170
rect 264 155 273 668
rect 363 629 372 668
rect 462 629 471 668
rect 363 195 372 580
rect 334 186 372 195
rect 334 155 343 163
rect 462 156 471 580
rect 528 428 537 668
rect 651 542 660 758
rect 689 683 698 758
rect 729 683 738 818
rect 767 807 776 818
rect 805 807 814 818
rect 767 746 776 758
rect 767 683 776 725
rect 805 683 814 758
rect 843 716 852 818
rect 881 807 890 818
rect 921 807 930 818
rect 881 746 890 783
rect 843 683 852 695
rect 881 683 890 725
rect 921 716 930 783
rect 921 683 930 695
rect 528 156 537 401
rect 651 311 660 521
rect 689 374 698 634
rect 729 598 738 634
rect 767 598 776 634
rect 805 598 814 634
rect 843 598 852 634
rect 729 513 738 549
rect 689 353 695 374
rect 651 231 660 290
rect 651 222 662 231
rect 653 210 662 222
rect 689 210 698 353
rect 729 317 738 492
rect 767 317 776 549
rect 805 350 814 549
rect 805 317 814 329
rect 843 317 852 549
rect 881 422 890 634
rect 921 422 930 634
rect 961 598 970 818
rect 961 479 970 549
rect 881 401 892 422
rect 881 317 890 401
rect 921 311 930 401
rect 653 170 662 183
rect 651 161 662 170
rect 66 59 75 128
rect 132 61 141 128
rect 198 63 207 128
rect 264 86 273 128
rect 334 88 343 128
rect 462 86 471 129
rect 528 65 537 129
rect 334 45 343 61
rect 651 48 660 161
rect 689 108 698 183
rect 729 141 738 290
rect 767 210 776 290
rect 805 210 814 290
rect 767 171 776 183
rect 729 108 738 120
rect 767 108 776 150
rect 805 108 814 183
rect 843 168 852 290
rect 881 204 890 290
rect 921 210 930 290
rect 843 108 852 144
rect 881 168 890 183
rect 921 168 930 183
rect 689 48 698 81
rect 729 48 738 81
rect 767 48 776 81
rect 805 48 814 81
rect 843 48 852 81
rect 881 48 890 144
rect 921 117 930 144
rect 961 117 970 458
rect 903 108 930 117
rect 943 108 970 117
rect 903 48 912 108
rect 943 93 952 108
rect 943 48 952 66
<< ndiffusion >>
rect 116 169 132 196
rect 141 169 146 196
rect 724 290 729 317
rect 738 290 767 317
rect 776 290 805 317
rect 814 290 817 317
rect 838 290 843 317
rect 852 290 881 317
rect 890 290 895 317
rect 650 183 653 210
rect 662 183 689 210
rect 698 183 703 210
rect 61 128 66 155
rect 75 128 132 155
rect 141 128 156 155
rect 177 128 198 155
rect 207 128 227 155
rect 250 128 264 155
rect 273 128 334 155
rect 343 128 386 155
rect 449 129 462 156
rect 471 129 528 156
rect 537 129 541 156
rect 328 61 334 88
rect 343 61 352 88
rect 764 183 767 210
rect 776 183 805 210
rect 814 183 817 210
rect 916 183 921 210
rect 930 183 935 210
rect 686 81 689 108
rect 698 81 729 108
rect 738 81 767 108
rect 776 81 805 108
rect 814 81 817 108
rect 838 81 843 108
rect 852 81 855 108
rect 938 66 943 93
rect 952 66 955 93
<< pdiffusion >>
rect 115 757 132 806
rect 141 757 160 806
rect 648 758 651 807
rect 660 758 665 807
rect 686 758 689 807
rect 698 758 703 807
rect 60 668 66 717
rect 75 668 93 717
rect 114 668 132 717
rect 141 668 161 717
rect 182 668 198 717
rect 207 668 226 717
rect 247 668 264 717
rect 273 668 323 717
rect 344 668 363 717
rect 372 668 381 717
rect 449 668 462 717
rect 471 668 490 717
rect 511 668 528 717
rect 537 668 541 717
rect 351 580 363 629
rect 372 580 387 629
rect 764 758 767 807
rect 776 758 781 807
rect 802 758 805 807
rect 814 758 817 807
rect 686 634 689 683
rect 698 634 703 683
rect 724 634 729 683
rect 738 634 743 683
rect 764 634 767 683
rect 776 634 781 683
rect 802 634 805 683
rect 814 634 817 683
rect 838 634 843 683
rect 852 634 855 683
rect 876 634 881 683
rect 890 634 895 683
rect 916 634 921 683
rect 930 634 935 683
rect 724 549 729 598
rect 738 549 743 598
rect 764 549 767 598
rect 776 549 781 598
rect 802 549 805 598
rect 814 549 817 598
rect 838 549 843 598
rect 852 549 855 598
rect 956 549 961 598
rect 970 549 973 598
<< pohmic >>
rect 0 30 603 32
rect 0 9 86 30
rect 107 9 157 30
rect 178 9 386 30
rect 409 9 456 30
rect 479 11 603 30
rect 624 11 1023 32
rect 479 9 1023 11
rect 0 7 1023 9
<< nohmic >>
rect 0 858 1023 859
rect 0 837 83 858
rect 104 837 155 858
rect 176 857 471 858
rect 176 837 406 857
rect 0 836 406 837
rect 429 837 471 857
rect 494 855 1023 858
rect 494 837 603 855
rect 429 836 603 837
rect 0 834 603 836
rect 624 834 1023 855
<< ntransistor >>
rect 132 169 141 196
rect 729 290 738 317
rect 767 290 776 317
rect 805 290 814 317
rect 843 290 852 317
rect 881 290 890 317
rect 653 183 662 210
rect 689 183 698 210
rect 66 128 75 155
rect 132 128 141 155
rect 198 128 207 155
rect 264 128 273 155
rect 334 128 343 155
rect 462 129 471 156
rect 528 129 537 156
rect 334 61 343 88
rect 767 183 776 210
rect 805 183 814 210
rect 921 183 930 210
rect 689 81 698 108
rect 729 81 738 108
rect 767 81 776 108
rect 805 81 814 108
rect 843 81 852 108
rect 943 66 952 93
<< ptransistor >>
rect 132 757 141 806
rect 651 758 660 807
rect 689 758 698 807
rect 66 668 75 717
rect 132 668 141 717
rect 198 668 207 717
rect 264 668 273 717
rect 363 668 372 717
rect 462 668 471 717
rect 528 668 537 717
rect 363 580 372 629
rect 767 758 776 807
rect 805 758 814 807
rect 689 634 698 683
rect 729 634 738 683
rect 767 634 776 683
rect 805 634 814 683
rect 843 634 852 683
rect 881 634 890 683
rect 921 634 930 683
rect 729 549 738 598
rect 767 549 776 598
rect 805 549 814 598
rect 843 549 852 598
rect 961 549 970 598
<< polycontact >>
rect 192 757 213 806
rect 326 792 347 818
rect 259 749 280 774
rect 60 401 81 426
rect 126 377 149 401
rect 191 170 213 194
rect 455 580 476 629
rect 322 163 346 186
rect 757 725 778 746
rect 881 783 905 807
rect 921 783 945 807
rect 873 725 894 746
rect 831 695 852 716
rect 909 695 930 716
rect 645 521 666 542
rect 519 401 545 428
rect 717 492 738 513
rect 695 353 716 374
rect 645 290 666 311
rect 800 329 821 350
rect 961 458 982 479
rect 916 401 937 422
rect 921 290 942 311
rect 256 65 281 86
rect 456 61 480 86
rect 757 150 778 171
rect 723 120 744 141
rect 869 183 890 204
rect 828 144 852 168
rect 881 144 905 168
rect 921 144 945 168
<< ndiffcontact >>
rect 95 169 116 196
rect 146 169 167 196
rect 703 290 724 317
rect 817 290 838 317
rect 895 290 916 317
rect 629 183 650 210
rect 703 183 724 210
rect 40 128 61 155
rect 156 128 177 155
rect 227 128 250 155
rect 386 128 407 155
rect 428 129 449 156
rect 541 129 562 156
rect 307 61 328 88
rect 352 61 373 88
rect 743 183 764 210
rect 817 183 838 210
rect 895 183 916 210
rect 935 183 956 210
rect 665 81 686 108
rect 817 81 838 108
rect 855 81 876 108
rect 917 66 938 93
rect 955 66 976 93
<< pdiffcontact >>
rect 94 757 115 806
rect 160 757 181 806
rect 627 758 648 807
rect 665 758 686 807
rect 703 758 724 807
rect 39 668 60 717
rect 93 668 114 717
rect 161 668 182 717
rect 226 668 247 717
rect 323 668 344 717
rect 381 668 402 717
rect 428 668 449 717
rect 490 668 511 717
rect 541 668 562 717
rect 330 580 351 629
rect 387 580 408 629
rect 743 758 764 807
rect 781 758 802 807
rect 817 758 838 807
rect 665 634 686 683
rect 703 634 724 683
rect 743 634 764 683
rect 781 634 802 683
rect 817 634 838 683
rect 855 634 876 683
rect 895 634 916 683
rect 935 634 956 683
rect 703 549 724 598
rect 743 549 764 598
rect 781 549 802 598
rect 817 549 838 598
rect 855 549 876 598
rect 935 549 956 598
rect 973 549 994 598
<< psubstratetap >>
rect 86 9 107 30
rect 157 9 178 30
rect 386 9 409 30
rect 456 9 479 30
rect 603 11 624 32
<< nsubstratetap >>
rect 83 837 104 858
rect 155 837 176 858
rect 406 836 429 857
rect 471 837 494 858
rect 603 834 624 855
<< metal1 >>
rect 0 858 1023 859
rect 0 837 83 858
rect 104 837 155 858
rect 176 857 471 858
rect 176 837 406 857
rect 0 836 406 837
rect 429 837 471 857
rect 494 855 1023 858
rect 494 837 603 855
rect 429 836 603 837
rect 0 834 603 836
rect 624 834 1023 855
rect 99 806 111 834
rect 181 757 192 806
rect 43 733 177 745
rect 43 717 55 733
rect 165 717 177 733
rect 230 717 242 834
rect 165 568 177 668
rect 299 608 311 834
rect 385 717 397 834
rect 627 807 639 834
rect 708 807 720 834
rect 748 807 760 834
rect 822 807 834 834
rect 433 737 557 749
rect 433 717 445 737
rect 545 717 557 737
rect 327 655 339 668
rect 495 655 507 668
rect 327 643 507 655
rect 299 596 330 608
rect 408 595 455 607
rect 545 568 557 668
rect 627 622 639 758
rect 669 740 681 758
rect 669 728 757 740
rect 790 740 802 758
rect 790 728 873 740
rect 894 728 956 740
rect 708 701 831 713
rect 708 683 720 701
rect 786 683 798 701
rect 864 701 909 713
rect 864 683 876 701
rect 944 683 956 728
rect 669 622 681 634
rect 748 622 760 634
rect 821 622 833 634
rect 899 622 911 634
rect 627 610 989 622
rect 748 598 760 610
rect 821 598 833 610
rect 977 598 989 610
rect 165 556 557 568
rect 876 586 935 598
rect 708 537 720 549
rect 786 537 798 549
rect 666 525 798 537
rect 176 499 567 511
rect 555 482 567 499
rect 860 509 872 549
rect 738 497 872 509
rect 555 470 674 482
rect 30 458 167 468
rect 662 458 961 470
rect 30 456 572 458
rect 30 446 42 456
rect 155 446 572 456
rect 0 434 42 446
rect 560 434 1023 446
rect 0 401 60 413
rect 647 413 893 422
rect 545 410 916 413
rect 545 401 659 410
rect 881 401 916 410
rect 937 401 1023 413
rect 0 377 126 389
rect 671 389 869 398
rect 149 386 1023 389
rect 149 377 683 386
rect 857 377 1023 386
rect 0 353 695 365
rect 716 365 845 374
rect 716 362 1023 365
rect 833 353 1023 362
rect 0 329 800 341
rect 821 329 1023 341
rect 666 290 703 302
rect 916 290 921 311
rect 821 256 833 290
rect 629 244 833 256
rect 96 220 108 232
rect 47 208 444 220
rect 47 155 59 208
rect 167 170 191 194
rect 99 32 111 169
rect 391 155 403 208
rect 432 156 444 208
rect 629 210 641 244
rect 743 210 755 244
rect 845 234 951 246
rect 845 222 857 234
rect 826 210 857 222
rect 939 210 951 234
rect 890 183 895 204
rect 161 32 173 128
rect 231 115 243 128
rect 544 115 556 129
rect 231 103 556 115
rect 373 67 456 79
rect 311 32 323 61
rect 629 32 641 183
rect 712 171 724 183
rect 712 159 757 171
rect 744 120 976 132
rect 670 108 682 120
rect 964 93 976 120
rect 876 81 917 93
rect 822 32 834 81
rect 0 30 603 32
rect 0 9 86 30
rect 107 9 157 30
rect 178 9 386 30
rect 409 9 456 30
rect 479 11 603 30
rect 624 11 1023 32
rect 479 9 1023 11
rect 0 7 1023 9
<< m2contact >>
rect 259 749 280 774
rect 93 674 114 700
rect 326 792 347 818
rect 881 783 905 807
rect 921 783 945 807
rect 154 495 176 519
rect 90 232 116 260
rect 322 163 346 186
rect 256 65 281 86
rect 828 144 852 168
rect 881 144 905 168
rect 921 144 945 168
rect 664 120 688 144
<< metal2 >>
rect 264 774 278 866
rect 330 818 344 866
rect 891 807 905 866
rect 924 807 938 866
rect 96 514 110 674
rect 96 500 154 514
rect 96 260 110 500
rect 891 168 905 783
rect 924 168 938 783
rect 264 0 278 65
rect 330 0 344 163
rect 688 130 852 144
rect 891 0 905 144
rect 924 0 938 144
<< labels >>
rlabel metal1 0 834 0 859 3 Vdd!
rlabel metal2 264 866 278 866 5 D
rlabel metal2 330 866 344 866 5 Load
rlabel metal2 330 0 344 0 1 Load
rlabel metal2 264 0 278 0 1 D
rlabel metal1 0 7 0 32 3 GND!
rlabel metal1 0 377 0 389 3 Test
rlabel metal1 0 353 0 365 3 Clock
rlabel metal1 0 329 0 341 3 nReset
rlabel metal1 0 401 0 413 3 SDI
rlabel metal1 0 434 0 446 3 ScanReturn
rlabel metal1 1023 434 1023 446 7 ScanReturn
rlabel metal1 1023 353 1023 365 7 Clock
rlabel metal1 1023 377 1023 389 7 Test
rlabel metal1 1023 401 1023 413 7 Q
rlabel metal1 1023 329 1023 341 7 nReset
rlabel metal1 1023 834 1023 859 7 Vdd!
rlabel metal1 1023 7 1023 32 7 GND!
rlabel metal2 891 0 905 0 1 nQ
rlabel metal2 924 0 938 0 1 Q
rlabel metal2 891 866 905 866 5 nQ
rlabel metal2 924 866 938 866 5 Q
<< end >>
